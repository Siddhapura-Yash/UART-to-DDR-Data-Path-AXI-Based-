module axi(
    //global signals
    input axi_clk,
    input rst,

    //extra internal signal
    input start,

    input [255:0] data_in,      //data will come from fifo
    input check_empty,          //empty signal from async fifo
    output read_enable,         //axi send read enable to the async fifo

    //Write address channel signals
    output [7:0] aid,           //transaction id
    output reg [31:0] aaddr,    //main address
    output reg [7:0] alen,      //burst length exact number of transfers (beats)
    output reg [2:0] asize,     //how wide each beat
    output reg [1:0] aburst,    //burst type(i.e fixed,wrap......)
    output reg [1:0] alock,     //00 for our case
    output reg avalid,          //valid signal master to slave 
    input aready,               //slave responds i'm ready to acccept addresss
    output reg atype,           //read or write 1 = write 0 = read

    // Write data channel signals
    output [7:0] wid,            //write transaction id
    output reg [255:0] wdata,    //actual write data
    output  [31:0] wstrb,        //write strobe
    output reg wlast,            //last data beat of burst
    output reg wvalid,           //high means write data is valid
    input wready,                //slave says i'm ready to accept data

    // Read data channel signals
    input [7:0] rid,            //read trasaction id
    input [255:0] rdata,        //read data from ddr
    input rlast,                //last beat of read burst
    input rvalid,               //high means read data is valid
    output reg rready,          //master ready to accepet read data
    input [1:0] rresp,          //read response 
									//00 → OKAY
									//01 → EXOKAY
									//10 → SLVERR
									//11 → DECERR

    // Write response channel signals                          
    input [7:0] bid,            //write response id
    input bvalid,               //Slave → Master high means write response is valid
    output reg bready,          //Master → Slave high means master ready to accept response 


    output reg fail,
    output reg done,
    output reg [255:0] obs_rdata_exp,
    output reg [255:0] obs_rdata_det,

    output [3:0]o_states
);

//will fetch data from word fifo
assign read_enable = !check_empty && wready;



assign aid = 8'h00;
assign wstrb = 32'hFFFFFFFF;
assign wid = 8'h00;

parameter ALEN = 23;
parameter ASIZE = 5;
parameter START_ADDR = 32'h00000000; 
parameter STOP_ADDR = 32'h00100000;
parameter ADDR_OFFSET = (ALEN + 1)*32;


//Main states
localparam
	IDLE = 4'b0000, 
	WRITE_ADDR = 4'b0001,
	PRE_WRITE = 4'b0010,
	WRITE = 4'b0011,
	POST_WRITE = 4'b0100,
	READ_ADDR = 4'b0101,
	PRE_READ = 4'b0110,
	READ_COMPARE = 4'b0111,
	POST_READ = 4'b1000,
	DONE = 4'b1001;

    reg [3:0] states, nstates;
    reg bvalid_done;
    reg [1:0] start_sync;
    reg [8:0] write_cnt, read_cnt;
    reg [255:0] rdata_store;
    reg wburst_done, rburst_done, write_done, read_done;

    always @(posedge axi_clk or negedge rstn) begin
        if (!rstn) begin
            start_sync <= 2'b00;
        end else begin
            start_sync[0] <= start;
            start_sync[1] <= start_sync[0];
        end
    end

    always @(posedge axi_clk or negedge rstn) begin
        if (!rstn) begin
        states <= IDLE;
        end else begin
        states <= nstates;
        end
    end

always @(states or start_sync[1] or write_cnt or rburst_done or write_done or read_done or bvalid_done or aready) begin
	case(states) 
	IDLE 	   : if (start_sync[1]) 			nstates = WRITE_ADDR;
	             else					nstates = IDLE;
	WRITE_ADDR : if (aready)				nstates = PRE_WRITE;
		     else					nstates = WRITE_ADDR;
	PRE_WRITE  : 						nstates = WRITE;
	WRITE	   : if (write_cnt == 9'd0)			nstates = POST_WRITE;
		     else		 			nstates = WRITE;
	POST_WRITE : if (write_done & bvalid_done) 		nstates = READ_ADDR;
		     else if (bvalid_done)			nstates = WRITE_ADDR;
		     else					nstates = POST_WRITE;
	READ_ADDR  : if (aready) 				nstates = PRE_READ;
		     else					nstates = READ_ADDR;
	PRE_READ   :						nstates = READ_COMPARE;
	READ_COMPARE  : if (rburst_done) 			nstates = POST_READ;
			else					nstates = READ_COMPARE;
	POST_READ  :	if (read_done) 				nstates = DONE;
			else					nstates = READ_ADDR;
	DONE	   : 						nstates = DONE;
	default							nstates = IDLE;
	endcase
end




always @(posedge axi_clk or negedge rstn) begin
	if (!rstn) begin
		aaddr <= START_ADDR;
		avalid <= 1'b0;
		atype <= 1'b0;
		aburst <= 2'b00;
		asize <= 3'b000;
		alen <= 8'd0;
		alock <= 2'b00;
		wvalid <= 1'b0;
		write_cnt <= ALEN + 1;
		write_done <= 1'b0;
		wdata <= 256'd0;
		wburst_done <= 1'b0;
		wlast <= 1'b0;
		bready <= 1'b0;
		fail <= 1'b0;
		done <= 1'b0;
		rready <= 1'b0;
		bvalid_done <=1'b0;
		obs_rdata_det <= 256'h0;
		obs_rdata_exp <= 256'h0;
	end else begin
		if (states == IDLE) begin
	                aaddr <= START_ADDR;
	                avalid <= 1'b0;
        	        atype <= 1'b0;
               	 	aburst <= 2'b00;
                	asize <= 3'b000;
                	alen <= 8'd0;
                	alock <= 2'b00;
                	wvalid <= 1'b0;
                	write_cnt <= ALEN + 1;
                	wdata <= 256'd0;
                	wburst_done <= 1'b0;
                	wlast <= 1'b0;
                	bready <= 1'b0;
			rready <= 1'b0;
			bvalid_done <= 1'b0;
			fail <= 1'b0;
			done <= 1'b0;
		end
		if (states == WRITE_ADDR) begin
			avalid <= 1'b1;
			atype <= 1'b1;
			asize <= ASIZE;
			alen <= ALEN;
			aburst <= 2'b01;
			alock <= 2'b00;
			wvalid <= 1'b0;
			write_cnt <= ALEN + 1;
			wburst_done <= 1'b0;
			bvalid_done <= 1'b0;
			bready <= 1'b0;
			rready <= 1'b0;
			done <= 1'b0;
			fail <= 1'b0;
		end
		if (states == PRE_WRITE) begin
			avalid <= 1'b0;
			atype <= 1'b0;
			wvalid <= 1'b1;
			wdata <= data_in;
			bready <= 1'b1;
			write_cnt <= write_cnt - 1;
            end
        if (states == WRITE) begin
                if (wready == 1'b1 && ) begin
                    wdata <= data_in;
                    if (write_cnt == 9'd0) begin
                    wburst_done <= 1'b1;
                    wlast <= 1'b0;
                    wvalid <= 1'b0;
                        if (aaddr >= STOP_ADDR) begin
                        write_done <= 1'b1;
                        end else begin
                        write_done <= 1'b0;
                        end
                    end if (write_cnt == 9'd1) begin
                        wlast <= 1'b1;
                        write_cnt <= write_cnt - 1;
                    end else begin
                    write_cnt <= write_cnt - 1;
                    end
                end
            end
            if (states == POST_WRITE) begin
                if (write_done) begin
                    aaddr <= START_ADDR;
                end else begin
                    if (bvalid) begin
                    aaddr <= aaddr + ADDR_OFFSET;
                    end
                end
                if (wready == 1'b1) begin
                    wlast <= 1'b0;	
                    wvalid <= 1'b0;	
                end
                if (bvalid) begin
                    bvalid_done <= 1'b1;
                    bready <= 1'b0;
                end
            end
            if (states == READ_ADDR) begin
                avalid <= 1'b1;
                read_cnt <= ALEN + 1;
                    
            end
            if (states == PRE_READ) begin
                avalid <= 1'b0;
                rburst_done <= 1'b0;
                            rdata_store <= {aaddr, ~aaddr, {8{~read_cnt[7:0]}},~aaddr,aaddr,{8{read_cnt[7:0]}}};
                read_cnt <= read_cnt - 1'b1;
            end
            if (states == READ_COMPARE) begin
                rready <= 1'b1;
                if (read_cnt != 9'd0) begin
                if (rvalid == 1'b1) begin
                            rdata_store <= {aaddr, ~aaddr, {8{~read_cnt[7:0]}},~aaddr,aaddr,{8{read_cnt[7:0]}}};
                read_cnt <= read_cnt - 1'b1;
                    if (rdata != rdata_store) begin
                        fail <= 1'b1;
                        obs_rdata_exp <= rdata_store;
                        obs_rdata_det <= rdata;
                        `ifdef EFX_SIM
                        $display("ERROR!! Read mismatch : read = 0x%x, expected = 0x%x",rdata,rdata_store);
                        `endif 
                    end else begin
                        `ifdef EFX_SIM
                        $display("Read match: read = 0x%x, expected = 0x%x",rdata,rdata_store);
                        `endif
                    end
        
                end
                end
                if (read_cnt == 9'd0) begin
                                if (rvalid == 1'b1) begin
                                        if (rdata != rdata_store) begin
                                                    fail <= 1'b1;

                                                    obs_rdata_exp <= rdata_store;

                                                    obs_rdata_det <= rdata;
                                                    `ifdef EFX_SIM
                                                    $display("ERROR!! Read mismatch : read = 0x%x, expected = 0x%x",rdata,rdata_store);
                                                    `endif
                                            end else begin
                                                    `ifdef EFX_SIM
                                                    $display("Read match: read = 0x%x, expected = 0x%x",rdata,rdata_store);
                                                    `endif
                                            end


                        if (aaddr >= STOP_ADDR) begin
                            read_done <= 1'b1;
                        end else begin
                            read_done <= 1'b0;
                        end
                        rburst_done <= 1'b1;
                    end
                end	
            end
            if (states == POST_READ) begin
                aaddr <= aaddr + ADDR_OFFSET;
                rready <= 1'b1;
            end
            if (states == DONE) begin
                done <= 1'b1;
            end
        end

    end


    assign o_states = states;

    endmodule